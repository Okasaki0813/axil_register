// SPDX-License-Identifier: CERN-OHL-S-2.0
/*

Copyright (c) 2018-2025 FPGA Ninja, LLC

Authors:
- Alex Forencich

*/

`resetall // ���ñ�������״̬��
          // Ϊʲô֮ǰ���ļ��ж���ĺ���ܻ�Ӱ�쵽��ǰ�ļ��ı��룿
          // �궨��ĳ�����ȫ�ֵ�
`timescale 1ns / 1ps
`default_nettype none // Ҫ�������źŶ�Ҫ��������ʹ�ã������������ֱ�ӱ���

/*
 * AXI4 lite register
 * ��ģ��������AXI-Lite�����ͨ����������Ĵ������ж�����߼�·��
 * ΪʲôҪ�üĴ����ж�����߼�·����������߼��������źſ����޷���һ��ʱ���������ܵ��յ㣬�Ӷ����ʱ��Υ��
 * �Ĵ���������ж�����߼�·���ģ���һ������߼������Ϊ����
 */
module taxi_axil_register #
(
    // 0 to bypass, 1 for simple buffer
    // 0��Bypass����·�������ģ�ֱ��͸��
    // ��1�ľ����ӳ�һ��ʱ������
    // ͸�������źŲ������κμĴ�����ֱ�Ӵ�����˵��������
    // 1��Simple buffer���򵥻���
    // Ϊʲô����һ��ʱ�����ڵ��ӳ������ڽ��͸�·�����߼�ѹ�����ӳ�����߼���
    // AW channel register type
    parameter AW_REG_TYPE = 1, // д��ַͨ���Ĵ�������
    // W channel register type
    parameter W_REG_TYPE = 1, // д����ͨ���Ĵ�������
    // B channel register type
    parameter B_REG_TYPE = 1, // д��Ӧͨ���Ĵ�������
    // AR channel register type
    parameter AR_REG_TYPE = 1, // ����ַͨ���Ĵ�������
    // R channel register type
    parameter R_REG_TYPE = 1 // ������ͨ���Ĵ�������
)
(
    input  wire logic    clk, // ȫ��ʱ���ź�
    input  wire logic    rst, // ȫ�ָ�λ�ź�

    /*
     * AXI4-Lite slave interface
     * �������������Ĵӻ��ӿڣ��������ǽ�������Master��ԭʼ����
     * ԭʼ������ָ��Master�����ġ�δ���κδ���������ġ�Э��ת����λ������ȣ����ź�
     * ��ԭʼ�������ָ�����Ĵ���ģ�鴦�����źţ�����ʱ�����
     */
    taxi_axil_if.wr_slv  s_axil_wr, // дͨ���ӻ���
    taxi_axil_if.rd_slv  s_axil_rd, // ��ͨ���ӻ���

    /*
     * AXI4-Lite master interface
     * ��������ӻ��������ӿڣ������ǽ����ĺ������ת����������Slave�������ڴ�����裨��ô֮ǰ�ᵽ��slave��ʲô�أ���
     */
    taxi_axil_if.wr_mst  m_axil_wr, // дͨ��������
    taxi_axil_if.rd_mst  m_axil_rd // ��ͨ��������
);

/*
 * ʵ����дͨ��������ģ��
 * ��ģ�鸺��AW��W��B����ͨ���ļĴ��߼�
 */
taxi_axil_register_wr #(
    .AW_REG_TYPE(AW_REG_TYPE),
    .W_REG_TYPE(W_REG_TYPE),
    .B_REG_TYPE(B_REG_TYPE)
)
axil_register_wr_inst (
    .clk(clk),
    .rst(rst),

    /*
     * AXI4-Lite slave interface
     */
    .s_axil_wr(s_axil_wr), // ���Ӵӻ���д�ӿ�

    /*
     * AXI4-Lite master interface
     */
    .m_axil_wr(m_axil_wr) // ����������д�ӿ�
);

/*
 * ʵ������ͨ��������ģ��
 * ��ģ�鸺��AR��R����ͨ���ļĴ��߼�
 */
taxi_axil_register_rd #(
    .AR_REG_TYPE(AR_REG_TYPE),
    .R_REG_TYPE(R_REG_TYPE)
)
axil_register_rd_inst (
    .clk(clk),
    .rst(rst),

    /*
     * AXI4-Lite slave interface
     */
    .s_axil_rd(s_axil_rd), // ���Ӵӻ�����ӿ�

    /*
     * AXI4-Lite master interface
     */
    .m_axil_rd(m_axil_rd) // ������������ӿ�
);

endmodule

`resetall
