`ifndef UVM_TEST_AXIL_REGISTER_BASE_TEST_SV
`define UVM_TEST_AXIL_REGISTER_BASE_TEST_SV

`include "uvm_macros.svh"

class axil_register_base_test extends uvm_test;
    `uvm_component_utils(axil_register_base_test)

    axil_register_env env;
    axil_register_config cfg; // ʵ�������ö���cfg

    // ��� parent ����Ĭ��ֵΪ null���������ԣ��������ʱ���봫 parent
    function new(string name = "axil_register_base_test", uvm_component parent = null);
        super.new(name, parent);
    endfunction

    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);

        // cfg �������������пռ�飬��ֹʹ�ÿվ�����������Ų�Ĵ���
        cfg = axil_register_config::type_id::create("cfg");
        if (cfg == null) begin
            `uvm_fatal("CFG_CREATE_FAIL", "Failed to create axil_register_config object!")
        end

        // ���cfg�Ƿ��top��ȡ��vif���������cfg������
        if(!uvm_config_db#(virtual taxi_axil_if)::get(this, "", "vif", cfg.vif)) begin
            `uvm_fatal("NOVIF", "Test layer cannot get virtual interface vif from config_db!")
        end else begin
            // ��������Ϣ���ɹ���ȡ vif ʱ��ӡȷ�ϣ����ڷ�����־׷�ٺ͵���
            `uvm_info("VIF_GET_SUCCESS", "Virtual interface vif acquired successfully from config_db!", UVM_MEDIUM)
        end

        // ʹ�� "env*" ȷ�� env ����������������� agent������ͨ��ͨ����õ�����
        uvm_config_db#(axil_register_config)::set(this, "env*", "cfg", cfg);

        env = axil_register_env::type_id::create("env", this);
    endfunction

    task run_phase(uvm_phase phase);
        super.run_phase(phase);
        // �������գ�����ļ��������� smoke_test ������ʵ��
    endtask

    // virtual function void end_of_elaboration_phase(uvm_phase phase);
    //        super.end_of_elaboration_phase(phase);
    //        uvm_top.print_topology(); // ��ӡuvm��֤�����Ĳ㼶�ṹ
    // endfunction
endclass

`endif // UVM_TEST_AXIL_REGISTER_BASE_TEST_SV