`ifndef AXIL_REGISTER_SCOREBOARD_SV
`define AXIL_REGISTER_SCOREBOARD_SV

`include "uvm_macros.svh"

class axil_register_scoreboard extends uvm_scoreboard;
    `uvm_component_utils(axil_register_scoreboard)

    int check_count;
    int error_count;

    axil_register_config cfg;

    uvm_tlm_analysis_fifo #(axil_register_transaction) exp_fifo; // uvm_tlm_analysis_fifo��һ�������湦�ܵ�����
                                                                 // #(axil_register_transaction)��ָ������Ҫ���ܵı�������
    uvm_tlm_analysis_fifo #(axil_register_transaction) act_fifo;

    function new(string name = "axil_register_scoreboard", uvm_component parent);
        super.new(name, parent);
    endfunction

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        exp_fifo = new("exp_fifo", this);
        act_fifo = new("act_fifo", this);
        
        if(!uvm_config_db#(axil_register_config)::get(this, "", "cfg", cfg)) begin
            `uvm_fatal("NOCFG", "Scoreboard cannot get configuration object from config_db!")
        end
    endfunction

    // ��run_phase�в��ϱȶ����������е�����
    virtual task run_phase(uvm_phase phase);
        axil_register_transaction exp_tr, act_tr;
        forever begin
            exp_fifo.get(exp_tr); // get������������õĺ����������Ǵ������л�ȡ����
            act_fifo.get(act_tr);

            if (exp_tr.compare(act_tr)) begin // compare�������ص���boolֵ��1������ͬ��0����ͬ
                `uvm_info("SCB", "Match! DUT sent what scoreboard received.", UVM_HIGH)
            end else begin
                `uvm_error("SCB", "Mismatch! Package corrupted at the DUT!")
            end
        end
    endtask
endclass

`endif // AXIL_REGISTER_SCOREBOARD_SV