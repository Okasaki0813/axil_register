class axil_register_write_seq extends uvm_sequence#(axil_register_transaction);
    `uvm_object_utils(axil_register_write_seq)

    // ��������������������� virtual sequence ��ʹ�� with Լ��
    rand bit [31:0] addr;
    rand bit [31:0] data;
    rand bit [3:0]  strb;

    function new(string name = "axil_register_write_seq");
        super.new(name);
    endfunction

    virtual task body();
        // ����һ�� transaction ����
        req = axil_register_transaction::type_id::create("req");
        
        start_item(req); // ��ʼ����
        
        // �������еı���ֵ���ݸ� transaction
        req.operation = axil_register_transaction::WRITE;
        req.addr      = this.addr;
        req.data      = this.data;
        req.strb      = this.strb;
        
        finish_item(req); // �������ֲ����͸� driver
    endtask
endclass