// adapter��RAL����������֮����ݷ���ٵĽ�ɫ
`ifndef AXIL_REGISTER_REG_ADAPTER_SV
`define AXIL_REGISTER_REG_ADAPTER_SV

`include "uvm_macros.svh"

class axil_register_reg_adapter extends uvm_reg_adapter;
    `uvm_object_utils(axil_register_reg_adapter);

    function new(string name = "axil_register_reg_adapter");    // ���function���ӷ���ֵ���ͣ�����ֵ��Ĭ��������1bit��logic
                                                                // ���ǹ��캯��������һ����������������������ֵ���ͣ���Ĭ�Ϸ��ظ���Ķ���ʵ��
        super.new(name);
        provides_responses = 0;
        supports_byte_enable = 1;
    endfunction

    // �� Sequence �е��� reg.write/read ʱ��UVM �Զ����ô˺���
    virtual function uvm_sequence_item reg2bus(const ref uvm_reg_bus_op rw); // const�ú����ڲ�ֻ�ܶ�ȡrw�����ݣ������޸���
                                                                             // ref��ʾ���ô���
                                                                             // uvm_reg_bus_op��uvm_reg���е�һ���ṹ��
                                                                             // ��uvm_reg_bus_op�Ķ�����ļ�ĩβ
                                                                            
        axil_register_transaction tr;
        tr = axil_register_transaction::type_id::create("tr");

        tr.operation = (rw.kind == UVM_WRITE) ? axil_register_transaction::WRITE : axil_register_transaction::READ;
        tr.addr      = rw.addr;
        tr.data      = rw.data;

        if (rw.kind == UVM_WRITE) begin
            tr.strb = rw.byte_en; // byte_en���ֽ�ʹ�ܣ����ڿ��ƼĴ������ʵ�����
        end else begin
            tr.strb = 4'b1111; // ������ʱ��д���������壬����Ϊȫ1
        end

        return tr;
    endfunction

    // ����������׽�����񲢷����� RAL ʱ��UVM �Զ����ô˺������¾���ֵ
    virtual function void bus2reg(uvm_sequence_item bus_item, ref uvm_reg_bus_op rw);
        axil_register_transaction tr;
        
        if(!$cast(tr, bus_item)) begin // cast����������ת������
            `uvm_fatal("ADAPT", $sformatf("bus_item type %s is not axil_register_transaction", 
                             bus_item.get_type_name()))
            return; // �˳���ǰ����
        end

        rw.kind    = (tr.operation == axil_register_transaction::WRITE) ? UVM_WRITE : UVM_READ;
        rw.addr    = tr.addr;
        rw.data    = tr.data;
        rw.byte_en = tr.strb;
        rw.status  = UVM_IS_OK;
    endfunction
endclass

`endif // AXIL_REGISTER_REG_ADAPTER_SV

// typedef struct {
//     uvm_access_e   kind;           // �������ͣ�UVM_READ �� UVM_WRITE
//     uvm_reg_addr_t addr;           // ��ַ��byte address��
//     uvm_reg_data_t data;           // ����
//     int            n_bits;         // �����ı�����
//     uvm_reg_byte_en_t byte_en;     // �ֽ�ʹ�ܣ�ÿ���ֽ�1bit��
//     uvm_status_e   status;         // ����״̬��UVM_IS_OK, UVM_HAS_X, UVM_NOT_OK
// } uvm_reg_bus_op;