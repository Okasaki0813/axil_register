`include "uvm_macros.svh"

class axil_register_monitor extends uvm_monitor;
    `uvm_component_utils(axil_register_monitor)

    virtual taxi_axil_if vif;

    uvm_analysis_port #(axil_register_transaction) ap; // �����˿����ڽ����ݰ���monitor������scoreboard

    function new(string name = "axil_register_monitor", uvm_component parent);
        super.new(name, parent);
        ap = new("ap", this);
    endfunction

    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);
    endfunction

    virtual task run_phase(uvm_phase phase);
        fork
            collect_write_data();
            collect_read_data();
        join
    endtask

    extern task collect_write_data();
    extern task collect_read_data();
endclass

task axil_register_monitor::collect_write_data();
    axil_register_transaction tr;

    forever begin
        tr = axil_register_transaction::type_id::create("tr"); // type_id��ʲô��create()������������ģ�
                                                               // type_id�ǹ����и����ֵ���ģ��
                                                               // create()�����պ��޸����еķ���ʱ�������Զ������µĶ��󣨹������ǣ�
        tr.operation = axil_register_transaction::WRITE;

        fork
            begin
                // ��׽д��ַAW
                wait(vif.awvalid === 1'b1 && vif.awready === 1'b1);
                tr.addr = vif.awaddr;
                tr.prot = vif.awprot;
                tr.user = vif.awuser;
            end

            begin
                // ��׽д����W
                wait(vif.wvalid === 1'b1 && vif.wready === 1'b1);
                tr.data = vif.wdata;
                tr.strb = vif.wstrb;
            end
        join

        // ��׽д��Ӧ
        wait(vif.bvalid === 1'b1 && vif.bready === 1'b1);
        tr.resp = vif.bresp;

        // �����ݷ��͸�scoreboard
        @(posedge vif.clk);
        ap.write(tr); // ���write������ap�Դ���
        `uvm_info(get_type_name(), "Collected a WRITE transaction", UVM_HIGH)
    end
endtask

task axil_register_monitor::collect_read_data();
    axil_register_transaction tr;

    forever begin
        tr = axil_register_transaction::type_id::create("tr");
        tr.operation = axil_register_transaction::READ;

        // ��׽����ַ�ź�AR
        wait(vif.arvalid === 1'b1 && vif.arready === 1'b1);
        tr.addr = vif.araddr;
        tr.prot = vif.arprot;
        tr.user = vif.aruser;

        // ��׽�������ź�R
        wait(vif.rvalid === 1'b1 && vif.rready === 1'b1);
        tr.data = vif.rdata;
        tr.resp = vif.rresp;

        @(posedge vif.clk);
        ap.write(tr);
    end
endtask