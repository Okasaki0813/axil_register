`ifndef AXIL_REGISTER_REG_BLOCK_SV
`define AXIL_REGISTER_REG_BLOCK_SV

`include "uvm_macros.svh"

class axil_register_reg_block extends uvm_reg_block;
    `uvm_object_utils(axil_register_reg_block)
    
    rand axil_register_reg_data  REG_DATA; // ʵ�����Ĵ���

    function new(string name = "axil_register_reg_block");
        super.new(name, UVM_NO_COVERAGE);
    endfunction

    virtual function void build();
        // �����Ĵ���ʵ��
        REG_DATA = axil_register_reg_data::type_id::create("REG_DATA");
        REG_DATA.configure(this, null, ""); // ���࣬����·��
        REG_DATA.build();

        // ������ַӳ��� (Address Map)
        // ���������֣�����ַ��ϵͳ����λ���ֽڣ����ֽ���
        default_map = create_map("default_map", 0, 4, UVM_LITTLE_ENDIAN);
        // ���Ĵ�������ӳ����Ĵ���ʵ����ƫ�Ƶ�ַ������Ȩ��
        default_map.add_reg(REG_DATA, 32'h0, "RW");
        
        lock_model(); // ����ģ�ͣ���ֹ��һ���޸�
    endfunction
endclass

`endif // AXIL_REGISTER_REG_BLOCK_SV