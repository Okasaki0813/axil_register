`include "uvm_macros.svh"

class axil_register_coverage extends uvm_subscriber #(axil_register_transaction);
    `uvm_component_utils(axil_register_coverage)

    axil_register_transaction m_item;
    
    covergroup axil_reg_cg; // ����������������ģ�Ϊʲôһ�������������ַ��˺ü���С�飿
        cp_operation: coverpoint m_item.operation { // m_item��ʲô������
            bins op_read  = {axil_register_transaction::READ};
            bins op_write = {axil_register_transaction::WRITE};
        }

        cp_addr: coverpoint m_item.addr { // ΪʲôҪ����ַ��Ϊ���ζ�����ֱ��һ���ж��ꣿ
            bins low_range    = {[32'h0000_0000 : 32'h0000_0FFF]};
            bins mid_range    = {[32'h0000_1000 : 32'hFFFF_EFFF]};
            bins high_range   = {[32'hFFFF_F000 : 32'hFFFF_FFFF]};
        }

        cp_strb: coverpoint m_item.strb { // Ϊʲôд����ֻ��ȫ1�Ͷ�������ʽ��������ʽ�أ�
            bins all_bytes = {4'b1111};
            bins single_byte = {4'b0001, 4'b0010, 4'b0100, 4'b1000};
        }

        cross_op_addr: cross cp_operation, cp_addr; // ʲô�ǽ��渲�ǣ�      
    endgroup

    function new(string name = "axil_register_coverage", uvm_component parent);
            super.new(name, parent);
            axil_reg_cg = new();
    endfunction  

    virtual function void write(axil_register_transaction t);
        m_item = t;
        axil_reg_cg.sample(); // ������ͨ����������ͳ�Ƹ�������
    endfunction
endclass