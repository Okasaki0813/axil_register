`include "uvm_macros.svh"

class axil_register_agent extends uvm_agent;
    `uvm_component_utils(axil_register_agent)

    virtual taxi_axil_if    vif;

    axil_register_sequencer sqr;
    axil_register_driver    drv;
    axil_register_monitor   mon;

    function new(string name = "axil_register_agent", uvm_component parent);
        super.new(name, parent);        
    endfunction

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);

        if(!uvm_config_db#(virtual taxi_axil_if)::get(this, "", "vif", vif)) begin  // get()�е��ĸ������ֱ���ʲô��˼��
                                                                                    // this�ǵ�ǰ�������monitor��ָ�룩
                                                                                    // ������Ѱ�Ҹ��ļ���ָ��·��
                                                                                    // ��vif����Ҫ�ҵ��ļ�������
                                                                                    // vif������ӿھ��
            `uvm_fatal("NOVIF", $sformatf("vif not found at path: %s", get_full_name()))
        end

        mon = axil_register_monitor::type_id::create("mon", this); // Ϊʲô�����create�������еڶ�������this�����Ǹ����õģ�
                                                                   // this����ָʾmon����ĸ�����������������uvm�Ĳ㼶�����ҵ���

        if(get_is_active() == UVM_ACTIVE) begin // get_is_active()��UVM_ACTIVE�ֱ���uvm_agent���õĺ����Ͳ������ǵ�
            sqr = axil_register_sequencer::type_id::create("sqr", this);
            drv = axil_register_driver::type_id::create("drv", this);
        end
    endfunction

    extern virtual function void connect_phase(uvm_phase phase); // Ϊʲô���������������ʵ�֣���Ҫ������ʵ�֣�
endclass

function void axil_register_agent::connect_phase(uvm_phase phase);
    super.connect_phase(phase);

    if (get_is_active() == UVM_ACTIVE) begin
        drv.vif = this.vif;
        drv.seq_item_port.connect(sqr.seq_item_export);
    end

    mon.vif = this.vif;
endfunction