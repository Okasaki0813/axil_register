`ifndef AXIL_REGISTER_TB_SV
`define AXIL_REGISTER_TB_SV

`include "uvm_macros.svh"

module axil_register_tb;
    logic clk;
    logic rst;

    // ����ʱ���źţ�Ƶ��Ϊ100MHz
    initial begin
        clk = 1'b0;
        forever #5 clk = ~clk;
    end

    // ���ɸ�λ�ź�
    // AXI4-Lite �и�λ�ǵ���Ч (active low)
    // rst = 1'b0: ��λ��Ч��ϵͳ���ڸ�λ״̬��
    // rst = 1'b1: ��λ�ͷţ�ϵͳ����������
    initial begin
        rst = 1'b0;      // ��ʼʱʩ�Ӹ�λ������Ч��
        #50 rst = 1'b1;  // �ȴ� 50ns ���ͷŸ�λ�������ֵĸ�λʱ���ַ������Ƿ���ַ����: ��ͬ��ַӳ����ȷ�ԡ�����/Խ���ַ����Ӧ��Ϊ��DECERR/SLVERR����
    end

    // Ϊ���� DUT �ڲ��� m_axil_* �� s_axil_* ���ӵ�ͬһ���ӿ�ʵ��
    //����ᵼ��ģ���ڲ���ͬһ�źŵ�˫������������ m_axil_wr.bready ��
    // ����ƽ̨������ bready ͬʱ����ͬһ net��������ʹ�������ӿ�ʵ����
    // - `master_if`�����ӵ� DUT ��������˿ڣ����� slave ��һ�ࣩ
    // - `slave_if` : ���ӵ� DUT �Ĵӻ���˿ڣ����� master ��һ�ࣩ
    // Testbench �� Master Agent Ӧʹ�� `slave_if`��Slave Agent ʹ�� `master_if`��
    taxi_axil_if #(
        .DATA_W(32),
        .ADDR_W(32)
    ) master_if(
        .clk(clk),
        .rst(rst)
    );

    taxi_axil_if #(
        .DATA_W(32),
        .ADDR_W(32)
    ) slave_if(
        .clk(clk),
        .rst(rst)
    );

    taxi_axil_register #(
        .AW_REG_TYPE(1),
        .W_REG_TYPE (1),
        .B_REG_TYPE (1),
        .AR_REG_TYPE(1),
        .R_REG_TYPE (1)
    ) dut (
        .clk(clk),
        .rst(rst),
        // ���ӣ�DUT �Ĵӻ��ڽӵ� `slave_if`��DUT �������ڽӵ� `master_if`
        .s_axil_wr(slave_if.wr_slv),
        .s_axil_rd(slave_if.rd_slv),
        .m_axil_wr(master_if.wr_mst),
        .m_axil_rd(master_if.rd_mst)
    );

    initial begin
        // Ϊ Test �����ýӿڣ�test ����Ҫ vif ����ȡ���ã�
        // ����ͬ�Ľӿ�ʵ���������ͬ�� agent��
        // - test �� Master Agent ʹ�� `slave_if`�������ӵ� DUT �Ĵӻ��ڣ���
        //   ��Ϊ Master Agent Ҫ�������� DUT ������s_axil_*����
        // - Slave Agent ʹ�� `master_if`�������ӵ� DUT �������ڣ���
        //   ��Ϊ Slave Agent ģ�����δ��豸������ m_axil_* �źš�
        uvm_config_db#(virtual taxi_axil_if)::set(null, "uvm_test_top*", "vif", slave_if);

        uvm_config_db#(virtual taxi_axil_if)::set(null, "uvm_test_top.env.agt*", "vif", slave_if);

        uvm_config_db#(virtual taxi_axil_if)::set(null, "uvm_test_top.env.slv_agt*", "vif", master_if);
        // null�������õ���ʼ·��
        // "uvm_test_top.env.slv_agt*"��Ŀ����������/����·��
        // vif����������ݿ��е�key
        // dut_if����Ҫ���ݵ�ʵ�ʶ�����

        run_test();
    end
endmodule

`endif // AXIL_REGISTER_TB_SV