`ifndef AXIL_SLAVE_DRIVER_SV
`define AXIL_SLAVE_DRIVER_SV

`include "uvm_macros.svh"

class axil_slave_driver extends axil_register_driver;
    `uvm_component_utils(axil_slave_driver)
    virtual taxi_axil_if vif; // ���鲻Ҫ�ڶ���ʱ�� modport���� connect ʱָ������

    function new(string name, uvm_component parent);
        super.new(name, parent);
    endfunction

    // ���� build_phase ����ȡ�ӿ�
    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase); // ������� super��ȷ������� get Ҳ��ִ�У�����еĻ���
        
        // �����ݿ��л�ȡ��Ϊ "vif" �Ľӿڣ�����ֵ�����ص� vif ����
        if (!uvm_config_db#(virtual taxi_axil_if)::get(this, "", "vif", vif)) begin
            `uvm_fatal("SLV_DRV", "Virtual interface not found for slave driver!")
        end
    endfunction
    
    // ��������������Ϊ Memory Model
    // ���ǵ�ַ��ֵ������
    bit [31:0] mem_model [bit [31:0]];

    virtual task run_phase(uvm_phase phase);
        bit aw_done = 1'b0; // д��ַͨ�����ֱ�־λ
        bit w_done  = 1'b0; // д����ͨ�����ֱ�־λ
        logic [31:0] saved_addr; // �����ݴ�awaddr����ֹ2��ʱ�����ں�vif.awaddr�����仯

        // ��ʼ����Slave Ĭ������ Ready
        vif.awready <= 1'b0;
        vif.wready  <= 1'b0;
        vif.bvalid  <= 1'b0;
        vif.arready <= 1'b0;
        vif.rvalid  <= 1'b0;

        forever begin
            @(posedge vif.clk);
            if (vif.rst) begin
                vif.bvalid  <= 1'b0;
                vif.awready <= 1'b0;
                vif.wready  <= 1'b0;
                vif.rvalid  <= 1'b0;
                aw_done     <= 1'b0;
                w_done      <= 1'b0;
            end else begin
                // Ĭ�ϱ��� Ready Ϊ 1 (ģ������ӻ�)
                vif.awready <= 1'b1;
                vif.wready  <= 1'b1;
                vif.arready <= 1'b1;

                // ģ�ⷴѹ��ÿ���� 30% �ĸ������� Ready��ģ��ӻ�æµ
                // vif.awready <= ( $urandom_range(0, 99) < 70 ); 
                // vif.wready  <= ( $urandom_range(0, 99) < 70 );
                // vif.arready <= ( $urandom_range(0, 99) < 70 );
                // `uvm_info("SLV_DRV", $sformatf("awready = 'b%0b, wready = 'b%0b, arready = 'b%0b", vif.awready, vif.wready, vif.arready), UVM_HIGH)
                
                // ע�⣺һ�� valid �� ready ���֣���һ��ͨ��Ҫ�����߼���
                // ����ļ���������ܵ������ֱ���������������Ҫ���Եġ�

                // ������׽��ͨ���������ź�
                if (vif.awvalid && vif.awready) begin 
                    aw_done = 1'b1;
                    saved_addr = vif.awaddr;
                end

                if (vif.wvalid && vif.wready)
                    w_done = 1'b1;

                // �����߼�����ַ�����ݶ����ֳɹ� (Valid & Ready ͬʱΪ 1)
                // if (vif.awvalid && vif.awready && vif.wvalid && vif.wready) begin   // ������ôд����Ϊд��ַ��д���ݺ�����ͬһ��ʱ�ӽ�����ͬʱ�������
                                                                                    // �������������д��ַͨ����д����ͨ�������ֳɹ��ź�        
                // `uvm_info("SLV_DRV", $sformatf("aw_done = 'b%0b, w_done = 'b%0b, vif.bvalid = 'b%0b", aw_done, w_done, vif.bvalid), UVM_HIGH)
                if (aw_done && w_done && !vif.bvalid) begin // ����!bvalid��Ϊ�˱�֤slave����Ӧ����master���ٴ�����һ������
                    // �ݴ浱ǰ��������ݣ���ֹ����һ�ĸ���
                    logic [31:0] addr_to_store = saved_addr;
                    logic [31:0] data_to_store = vif.wdata; // ��������ͨ����ʱ�ȶ�
                    logic [31:0] wstrb_mask;    // 32λ����
                    logic [31:0] old_data;      // ԭ������
                    logic [31:0] new_combined_data;

                    // �������״̬λ��׼��������һ������ 
                    aw_done = 1'b0; 
                    w_done  = 1'b0;

                    addr_to_store = saved_addr;

                    // ���� 32 λ���룺����λ���Ƽ���
                    // �� wstrb ��ÿһλ��չΪ 8 λ
                    wstrb_mask = {{8{vif.wstrb[3]}}, {8{vif.wstrb[2]}}, {8{vif.wstrb[1]}}, {8{vif.wstrb[0]}}};

                    // ��ȡ�����ݣ������������Ĭ��Ϊ0��
                    old_data = mem_model.exists(addr_to_store) ? mem_model[addr_to_store] : 32'h0;

                    // ������ݣ�(������ & ����) | (������ & ~����)
                    new_combined_data = (vif.wdata & wstrb_mask) | (old_data & ~wstrb_mask);

                    // ���´洢
                    mem_model[addr_to_store] = new_combined_data;

                    `uvm_info("SLV_MEM", $sformatf("WSTRB Write: Addr='h%0h, Data='h%0h, Mask='b%04b, Final='h%0h", 
                    addr_to_store, vif.wdata, vif.wstrb, new_combined_data), UVM_HIGH)

                    fork
                        begin
                            automatic logic [31:0] current_awaddr = saved_addr;
                            repeat(2) @(posedge vif.clk);   // ģ��ӻ��ӳ�
                                                            // ����ȴ����ܻᵼ��slave�޷���⵽master���͵��µ������źţ��Ӷ�©������
                                                            // ���������ʹ��fork-join_none�ṹ
                            vif.bvalid <= 1'b1;
                            vif.bresp  <= (current_awaddr > 32'h3FFF) ? 2'b10 : 2'b00;
                        
                            // ��Ӧ���ֳɹ���Master ���յ� (bready=1)��Slave ���� bvalid
                            do begin
                                @(posedge vif.clk);
                            end while (!vif.bready);

                            vif.bvalid <= 1'b0;
                        end
                    join_none
                end

                if (vif.arvalid && vif.arready && !vif.rvalid) begin;
                    `uvm_info("SLV_DRV", $sformatf("Read request received at addr 'h%0h", vif.araddr), UVM_LOW)

                    fork
                        begin
                            automatic logic [31:0] current_araddr = vif.araddr;
                            repeat(2) @(posedge vif.clk);
                            vif.rvalid <= 1'b1;
                            vif.rresp  <= (current_araddr > 32'h0000_3FFF) ? 2'b10 : 2'b00;                
                            // --- ��̬��ȡ�洢ģ�� ---
                            if (mem_model.exists(current_araddr)) begin
                                vif.rdata <= mem_model[current_araddr]; // ����֮ǰд����ֵ
                            end else begin
                                vif.rdata <= 32'hDEAD_BEEF; // ���ûд��������һ������ֵ��ʾ��δ���塱
                            end

                            do begin
                                @(posedge vif.clk);
                            end while(!vif.rready);

                            vif.rvalid <= 1'b0;
                        end
                    join_none
                end
            end
        end
    endtask
endclass

`endif // AXIL_SLAVE_DRIVER_SV