`ifndef AXIL_REGISTER_RESET_VIRT_SEQ_SV
`define AXIL_REGISTER_RESET_VIRT_SEQ_SV

`include "uvm_macros.svh"

// axil_register_reset_virt_seq.sv
// ��λ�������� - ����ʩ�Ӹ�λ�źŲ���֤ϵͳ��λ���״̬
class axil_register_reset_virt_seq extends axil_register_base_virtual_sequence;
    `uvm_object_utils(axil_register_reset_virt_seq)

    function new(string name = "axil_register_reset_virt_seq");
        super.new(name);
    endfunction

    virtual task body();
        int reset_cycles = 5;      // ��λ����ʱ�䣨ʱ����������
        int wait_after_reset = 10; // ��λ�ͷź�ĵȴ�ʱ��
        int cycle_cnt = 0;

        `uvm_info(get_type_name(), $sformatf("Starting Reset Sequence (reset for %0d cycles)...", reset_cycles), UVM_LOW)

        // ���� 1���ȴ���ʼ״̬�ȶ�����ѡ��ͨ������һ��ʼ���Ǹ�λ״̬��
        @(posedge p_sequencer.vif.clk);
        #1ps; // �ȴ� clock �������ȶ�

        // ���� 2���۲츴λ��ʩ�ӣ�rst �ɶ�������������ֻ�۲죩
        if (p_sequencer.vif.rst !== 1'b0) begin
            `uvm_warning(get_type_name(), "Expected rst=0 at start (topmodule should drive rst), but got rst=1")
        end

        // ���� 3���ȴ���λ�͵�ƽά��ָ����������
        `uvm_info(get_type_name(), $sformatf("Observing reset (low) for %0d clocks...", reset_cycles), UVM_LOW)
        repeat(reset_cycles) begin
            @(posedge p_sequencer.vif.clk);
            cycle_cnt++;
        end

        // ���� 4���ȴ���λ�źű��ͷţ��ɶ����ͷţ�
        `uvm_info(get_type_name(), "Waiting for reset to be released by topmodule...", UVM_LOW)
        wait(p_sequencer.vif.rst === 1'b1); // ����ֱ�� rst ���ͷ�
        @(posedge p_sequencer.vif.clk);
        #1ps; // �ȶ�

        // ���� 5���ȴ� N ������ʹϵͳ�ȶ�����
        `uvm_info(get_type_name(), $sformatf("Waiting %0d clocks for stabilization...", wait_after_reset), UVM_LOW)
        repeat(wait_after_reset) begin
            @(posedge p_sequencer.vif.clk);
        end

        // ���� 6����֤��λ���״̬
        `uvm_info(get_type_name(), "Verifying post-reset state...", UVM_LOW)
        verify_reset_state();

        `uvm_info(get_type_name(), "Reset Sequence PASSED", UVM_LOW)
    endtask

    // ��֤��������鸴λ�����������ź��Ƿ�ص���ʼ״̬
    virtual task verify_reset_state();
        bit pass = 1;

        // valid �ź�Ӧ��Ϊ 0������Ч����
        if (p_sequencer.vif.awvalid !== 1'b0) begin
            `uvm_error(get_type_name(), "awvalid signal not reset to 0")
            pass = 0;
        end
        if (p_sequencer.vif.wvalid !== 1'b0) begin
            `uvm_error(get_type_name(), "wvalid signal not reset to 0")
            pass = 0;
        end
        if (p_sequencer.vif.arvalid !== 1'b0) begin
            `uvm_error(get_type_name(), "arvalid signal not reset to 0")
            pass = 0;
        end

        // Ready signals can be any value (implementation dependent), but typically should be 0 or stable 1
        if (p_sequencer.vif.bvalid !== 1'b0) begin
            `uvm_warning(get_type_name(), "bvalid is not 0 (may be a design characteristic)")
        end
        if (p_sequencer.vif.rvalid !== 1'b0) begin
            `uvm_warning(get_type_name(), "rvalid is not 0 (may be a design characteristic)")
        end

        if (pass) begin
            `uvm_info(get_type_name(), "Post-reset state verification PASSED", UVM_LOW)
        end else begin
            `uvm_error(get_type_name(), "Post-reset state verification FAILED")
        end
    endtask

endclass

`endif // AXIL_REGISTER_RESET_VIRT_SEQ_SV