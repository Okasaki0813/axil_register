`ifndef AXIL_REGISTER_RAL_FIELD_VIRT_SEQ_SV
`define AXIL_REGISTER_RAL_FIELD_VIRT_SEQ_SV

class axil_register_ral_field_virt_seq extends axil_register_base_virtual_sequence;
    `uvm_object_utils(axil_register_ral_field_virt_seq)

    function new(string name = "axil_register_ral_field_virt_seq");
        super.new(name);
    endfunction

    virtual task body();
        uvm_status_e status;

        if (rm == null) `uvm_fatal("RAL_SEQ", "rm handle is null!")
        
        `uvm_info(get_type_name(), "Starting RAL Field-level Access Sequence...", UVM_LOW)

        // ���� 1: ͨ�� RAL ���Ĵ���дһ������ֵ (ȫ��д)
        // ��ʱ Adapter Ӧ���Զ����� strb = 4'b1111
        rm.REG_DATA.write(status, 32'h1122_3344, UVM_FRONTDOOR);

        // ���� 2: ���޸ļĴ����е�ĳ���ֶ� (Field-level update)
        // ��������Ҫ�ѵ� 16 λ�޸�Ϊ 0xAAAA
        // ע�⣺����ʹ�� set() ֻ�ı�ģ������ֵ�����������߶���
        rm.REG_DATA.fld_low.set(16'hAAAA);
        
        // ���� 3: ͬ��ģ�͵�Ӳ�� (update)
        // RAL ��ԱȾ���ֵ (h11223344) ������ֵ (hXXXXAAAA)
        // �����Զ�����ֻ�е������ֽڱ��ˣ��Ӷ�����һ������ strb = 4'b0011 �� AXI д����
        rm.REG_DATA.update(status);

        // ���� 4: ǰ�Ŷ�ȡ��֤
        rm.REG_DATA.mirror(status, UVM_CHECK, UVM_FRONTDOOR);
    endtask
endclass

`endif