`ifndef AXIL_REGISTER_RAL_FIELD_TEST_SV
`define AXIL_REGISTER_RAL_FIELD_TEST_SV

class axil_register_ral_field_test extends axil_register_base_test;
    `uvm_component_utils(axil_register_ral_field_test)

    function new(string name = "axil_register_ral_field_test", uvm_component parent);
        super.new(name, parent);
    endfunction

    // ��д run_phase��ʹ�� RAL ���ֶη��� API
    virtual task run_phase(uvm_phase phase);
        uvm_status_e status;
        uvm_reg_data_t data;

        phase.raise_objection(this);
        
        `uvm_info("FIELD_TEST", "Step 1: Write initial background value 32'h11223344", UVM_LOW)
        env.rm.REG_DATA.write(status, 32'h1122_3344, UVM_FRONTDOOR);

        // �ֶ���ģ��״̬��Ϊ����Ӳ��һ���Ҹɾ���
        env.rm.REG_DATA.predict(32'h1122_3344);

        `uvm_info("FIELD_TEST", "Step 2: Update only fld_low to 16'hAAAA", UVM_LOW)
        // ʹ�� set() ���ı�ģ���ڲ�����ֵ (Desired Value)
        env.rm.REG_DATA.fld_low.set(16'hAAAA);
        
        // ���� update()��RAL �ᷢ�� fld_high û�䣬ֻ�� fld_low ���� (Dirty)
        // ���� Adapter �� reg2bus ���յ�һ�� byte_en=4'b0011 ������
        env.rm.REG_DATA.update(status);

        #100ns;

        `uvm_info("FIELD_TEST", "Step 3: Mirror check. Expected Final Value: 32'h1122AAAA", UVM_LOW)
        env.rm.REG_DATA.mirror(status, UVM_CHECK, UVM_FRONTDOOR);

        phase.drop_objection(this);
    endtask
endclass

`endif