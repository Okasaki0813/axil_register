`ifndef AXIL_REGISTER_RESET_TEST_SV
`define AXIL_REGISTER_RESET_TEST_SV

// ��λ���� - ��֤ģ�鸴λ��ĳ�ʼ��״̬
class axil_register_reset_test extends axil_register_base_test;
    `uvm_component_utils(axil_register_reset_test)

    function new(string name = "axil_register_reset_test", uvm_component parent = null);
        super.new(name, parent);
    endfunction

    // ��ѡ���� build_phase ���Զ�������
    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        // ���ڴ˴����� scoreboard �� coverage��רע�ڸ�λ��֤
        // cfg.enable_scb = 0;
        // cfg.enable_cov = 0;
    endfunction

    // �������߼���������λ����
    virtual task run_phase(uvm_phase phase);
        axil_register_reset_virt_seq reset_seq = axil_register_reset_virt_seq::type_id::create("reset_seq");
        
        phase.raise_objection(this); // ���� UVM ����л���У���ֹ��ǰ��������
        
        `uvm_info(get_type_name(), "Starting Reset Test...", UVM_LOW)
        reset_seq.start(env.virt_sqr); // ������ sequencer ��ִ�и�λ����
        `uvm_info(get_type_name(), "Reset Test Completed", UVM_LOW)
        
        phase.drop_objection(this); // ���� UVM ��ܻ�ѽ���
    endtask

    // ��ѡ���� check_phase �н������յ���֤�͸�����ͳ��
    function void check_phase(uvm_phase phase);
        super.check_phase(phase);
        `uvm_info(get_type_name(), "Reset Test Check Phase - All verifications passed", UVM_LOW)
    endfunction

endclass

`endif // AXIL_REGISTER_RESET_TEST_SV
