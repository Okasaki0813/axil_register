class axil_register_random_test extends axil_register_base_test;
    `uvm_component_utils(axil_register_random_test)

    function new(string name = "axil_register_random_test", uvm_component parent); // test�ĸ������uvm_top
        super.new(name, parent);
    endfunction

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
    endfunction

    virtual task run_phase(uvm_phase phase);
        axil_register_random_virt_seq vseq = axil_register_random_virt_seq::type_id::create("vseq"); // create�����ǹ����ṩ�ģ��������Ǵ���һ������Ϊrandom_virt_seq������Ϊvseq��ʵ������
        phase.raise_objection(this);
        vseq.start(env.virt_sqr); // ���������˼������env�е�virt_sqr��ʼ�����������
        phase.drop_objection(this);
    endtask
endclass