class axil_register_base_virtual_sequence extends uvm_sequence;
    `uvm_object_utils(axil_register_base_virtual_sequence)

    axil_register_reg_block rm;
    
    `uvm_declare_p_sequencer(axil_register_virtual_sequencer) // �����������virtual sequence��Ȩ�޷���virtual sequencer�ڲ���agent

    function new(string name = "axil_register_base_virtual_sequence");
        super.new(name);
    endfunction

    // ����ͨ�����Է�һЩ���о籾ͨ�õĵȴ���λ��ɵ��߼�
    virtual task body();
        `uvm_info(get_type_name(), "Base virtual sequence body started", UVM_LOW)
    endtask
endclass