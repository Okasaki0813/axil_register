`include "uvm_macros.svh"

// axil_register_agent (deprecated)
// ���ݰ�װ: ����ԭ�� axil_register_agent �Ա��������/�ɴ�������ʧЧ��
// �Ƽ�ʹ�� `axil_register_master_agent`���˰�װ��̳��� `axil_register_master_agent` ������ԭĬ�����ơ�

class axil_register_agent extends axil_register_master_agent;
    `uvm_component_utils(axil_register_agent)

    function new(string name = "axil_register_agent", uvm_component parent = null);
        super.new(name, parent);
    endfunction
endclass