`ifndef AXIL_REGISTER_REG_PREDICTOR_SV
`define AXIL_REGISTER_REG_PREDICTOR_SV

`include "uvm_macros.svh"

// 1. �����Ҫ�İ�������������Ŀ������
import uvm_pkg::*;

// 2. ��������transaction�ࣨ��������axil_register_transaction��
`include "../../vip_lib/transactions/axil_register_transaction.sv"

// 3. ����adapter����Ϊpredictor��Ҫ��ͬ��adapter��
`include "axil_register_reg_adapter.sv"

class axil_register_reg_predictor extends uvm_reg_predictor#(axil_register_transaction);
    `uvm_component_utils(axil_register_reg_predictor)

    bit enable_prediction = 1; // �Ƿ�����Ԥ�⹦��
    bit debug_enable      = 0; // �Ƿ����õ������

    int num_predicted_writes = 0; // Ԥ���д��������
    int num_predicted_reads  = 0; // Ԥ��Ķ���������
    int num_predicted_errors = 0; // Ԥ��Ĵ�������

    function new(string name = "axil_register_reg_predictor", uvm_component parent = null);
        super.new(name, parent);
    endfunction

    virtual function void write(axil_register_transaction tr);
        if (!enable_prediction) begin
            `uvm_warning(get_type_name(), "Prediction is disabled, ignoring transaction")
            return;
        end

        super.write(tr); // ���ø����д��������Ԥ��

        if (tr.operation == axil_register_transaction::WRITE) begin
            num_predicted_writes++;
            if (debug_enable) begin
                `uvm_info(get_type_name(), 
                    $sformatf("Predicted WRITE: addr=0x%0h, data=0x%0h, strb=0x%0h", 
                    tr.addr, tr.data, tr.strb), 
                    UVM_HIGH)
            end
        end else begin
            num_predicted_reads++;
            if (debug_enable) begin
                `uvm_info(get_type_name(), 
                    $sformatf("Predicted READ: addr=0x%0h, data=0x%0h", 
                    tr.addr, tr.data), 
                    UVM_HIGH)
            end
        end
    endfunction
endclass

`endif // AXIL_REGISTER_REG_PREDICTOR_SV