// adapter��RAL����������֮����ݷ���ٵĽ�ɫ
`ifndef AXIL_REGISTER_REG_ADAPTER_SV
`define AXIL_REGISTER_REG_ADAPTER_SV

`include "uvm_macros.svh"

class axil_register_reg_adapter extends uvm_reg_adapter;
    `uvm_object_utils(axil_register_reg_adapter);

    function new(string name = "axil_register_reg_adapter");    // ���function���ӷ���ֵ���ͣ�����ֵ��Ĭ��������1bit��logic
                                                                // ���ǹ��캯��������һ����������������������ֵ���ͣ���Ĭ�Ϸ��ظ���Ķ���ʵ��
        super.new(name);
        provides_responses = 0;
        supports_byte_enable = 1;
    endfunction

    // �� Sequence �е��� reg.write/read ʱ��UVM �Զ����ô˺���
    virtual function uvm_sequence_item reg2bus(const ref uvm_reg_bus_op rw); // const�ú����ڲ�ֻ�ܶ�ȡrw�����ݣ������޸���
                                                                             // ref��ʾ���ô���
                                                                             // uvm_reg_bus_op��uvm_reg���е�һ���ṹ��
                                                                            
        axil_register_transaction tr;
        tr = axil_register_transaction::type_id::create("tr");

        tr.operation = (rw.kind == UVM_WRITE) ? axil_register_transaction::WRITE : axil_register_transaction::READ;
        tr.addr      = rw.addr;
        tr.data      = rw.data;

        if (rw.kind == UVM_WRITE) begin
            tr.strb = rw.byte_en;
        end else begin
            tr.strb = 4'b0000;
        end

        return tr;
    endfunction

    // ����������׽�����񲢷����� RAL ʱ��UVM �Զ����ô˺������¾���ֵ
    virtual function void bus2reg(uvm_sequence_item bus_item, ref uvm_reg_bus_op rw);
        axil_register_transaction tr;
        
        if(!$cast(tr, bus_item)) begin // cast����������ת������
            `uvm_fatal("ADAPT", "Provided bus_item is not of the correct type") // Ϊʲô���ﲻ��get_type_name�ˣ�
            return; // �˳���ǰ����
        end

        rw.kind   = (tr.operation == axil_register_transaction::WRITE) ? UVM_WRITE : UVM_READ;
        rw.addr   = tr.addr;
        rw.data   = tr.data;
        rw.status = UVM_IS_OK;
    endfunction
endclass

`endif // AXIL_REGISTER_REG_ADAPTER_SV