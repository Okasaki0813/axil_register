`ifndef AXIL_REGISTER_MASTER_AGENT_SV
`define AXIL_REGISTER_MASTER_AGENT_SV

`include "uvm_macros.svh"

// axil_register_master_agent
// ˵��: �������� axil_register_agent����Ϊ Master ��� UVM agent��
// ���ļ���ԭ�߼�һ�£��������Ա��� Slave/���� agent ���֡�
class axil_register_master_agent extends uvm_agent;
    `uvm_component_utils(axil_register_master_agent)

    // ����ӿھ������ testbench �� config_db ������
    virtual taxi_axil_if    vif;

    axil_register_sequencer sqr;
    axil_register_driver    drv;
    axil_register_monitor   mon;

    function new(string name = "axil_register_master_agent", uvm_component parent = null);
        super.new(name, parent);
    endfunction

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);

        // uvm_config_db::get(scope, inst_name, field_name, value)
        // - scope (this): �ӵ�ǰ�����ʼ��������
        // - inst_name (""): ���ַ�����ʾͨ�䣬���������Ӳ㼶
        // - field_name ("vif"): �� set ʱʹ�õļ�����Ӧ
        // - vif: ��������ӿھ���ı���
        if(!uvm_config_db#(virtual taxi_axil_if)::get(this, "", "vif", vif)) begin
            `uvm_fatal("NOVIF", $sformatf("vif not found at path: %s", get_full_name()))
        end

        // create(name, parent) �еĵڶ�����������ָ���������owner��
        // ������ҵ�������£����� UVM �㼶�������� reporting/configuration/path ��ѯ
        mon = axil_register_monitor::type_id::create("mon", this);

        // ���� agent ���ڼ���״̬��UVM_ACTIVE��ʱ���� sequencer �� driver
        if(get_is_active() == UVM_ACTIVE) begin
            sqr = axil_register_sequencer::type_id::create("sqr", this);
            drv = axil_register_driver::type_id::create("drv", this);
        end
    endfunction

    // ����������������������ʵ���� SystemVerilog/UE���÷��֮һ��
    // - �����ඨ���������
    // - ���ڰ�ʵ�ַ����ļ��ײ��򵥶��ļ���ʵ��
    extern virtual function void connect_phase(uvm_phase phase);
endclass

function void axil_register_master_agent::connect_phase(uvm_phase phase);
    super.connect_phase(phase);

    // ���� agent ����ʱ������ driver ������ӿ��� sequencer �Ķ˿�
    if (get_is_active() == UVM_ACTIVE) begin
        drv.vif = this.vif; // ���ӿھ�����ݸ� driver
        drv.seq_item_port.connect(sqr.seq_item_export); // ���� sequencer <-> driver
    end

    // monitor ������Ҫ�ӿ��Թ۲��źţ����ҲҪ���� vif
    mon.vif = this.vif;
endfunction

`endif // AXIL_REGISTER_MASTER_AGENT_SV
