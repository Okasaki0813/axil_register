// �Ĵ����Ĺ����������𽫶��uvm_regʵ����֯��һ�𣬲��������ǵĻ���ַ�͵�ַӳ���
`ifndef AXIL_REGISTER_REG_DATA_SV
`define AXIL_REGISTER_REG_DATA_SV

import uvm_pkg::*;
`include "uvm_macros.svh"

class axil_register_reg_data extends uvm_reg;
    `uvm_object_utils(axil_register_reg_data)

    rand uvm_reg_field fld_low;
    rand uvm_reg_field fld_high;

    function new(string name = "axil_register_reg_data");
        // ���������֣���λ���Ƿ�֧�ָ�����
        super.new(name, 32, UVM_NO_COVERAGE);
    endfunction

    virtual function void build();
        fld_low = uvm_reg_field::type_id::create("fld_low");
        // ���������࣬λ�����λλ�ã�����Ȩ�ޣ��Ƿ���ʧ����λֵ���Ƿ��и�λ���Ƿ��������Ƿ�ɵ�����ȡ
        fld_low.configure(this, 16, 0, "RW", 0, 16'h0, 1, 1, 1);

        fld_high = uvm_reg_field::type_id::create("fld_high");
        // ע�⣺��ʼλ����Ϊ 16
        fld_high.configure(this, 16, 16, "RW", 0, 16'h0, 1, 1, 1);
    endfunction
endclass

`endif // AXIL_REGISTER_REG_DATA_SV