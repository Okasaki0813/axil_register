class axil_register_smoke_virt_seq extends axil_register_base_virtual_sequence;
    // ð�̲�������֤��������򵥡�������Ĳ�������������Ҫ������֤����ͨ·
    `uvm_object_utils(axil_register_smoke_virt_seq)

    function new(string name = "axil_register_smoke_virt_seq");
        super.new(name);
    endfunction

    virtual task body();
        // ���������ײ��ԭ����������
        axil_register_write_seq  wr_seq;
        axil_register_read_seq   rd_seq;

        `uvm_info(get_type_name(), "Executing Smoke Virtual Sequence...", UVM_LOW)
        // get_type_name���ڻ�ȡ��������get_full_name���ڻ�ȡʵ����
        
        // 1. ִ��д����
        `uvm_do_on_with(wr_seq, p_sequencer.agt_sqr, {
            addr == 32'h0000_0004;
            data == 32'hAAAA_BBBB;
        })

        // 2. ִ�ж����������ղ�д�ĵ�ַ��
        `uvm_do_on_with(rd_seq, p_sequencer.agt_sqr, {
            addr == 32'h0000_0004;
        })
        
        `uvm_info(get_type_name(), "Smoke Virtual Sequence finished", UVM_LOW)
    endtask
endclass