`include "uvm_macros.svh"

// `include "taxi_axil_if.sv"
// `include "axil_register_transaction.sv"
// `include "axil_register_base_test.sv"

module top;
    logic clk;
    logic rst;

    // ����ʱ���źţ�Ƶ��Ϊ100MHz
    initial begin
        clk = 1'b0;
        forever #5 clk = ~clk;
    end

    // ���ɸ�λ�ź�
    initial begin
        rst = 1'b1;
        #20 rst = 1'b0;
    end

    taxi_axil_if #(
        .DATA_W(32),
        .ADDR_W(32)
    ) dut_if(
        .clk(clk),
        .rst(rst)
    );

    taxi_axil_register #(
        .AW_REG_TYPE(1),
        .W_REG_TYPE (1),
        .B_REG_TYPE (1),
        .AR_REG_TYPE(1),
        .R_REG_TYPE (1)
    ) dut (
        .clk(clk),
        .rst(rst),
        .s_axil_wr(dut_if.wr_slv),
        .s_axil_rd(dut_if.rd_slv),
        .m_axil_wr(dut_if.wr_mst),
        .m_axil_rd(dut_if.rd_mst)
    );

//     initial begin
//         uvm_config_db#(virtual taxi_axil_if)::set(null, "uvm_test_top.*", "vif", dut_if); // ���ĸ������ֱ���ʲô��˼��
//                                                                                           // null��������·��
//                                                                                           // uvm_test_top:*��Ŀ��·��
//                                                                                           // vif��key
//                                                                                           // dut_if��value
//         // �� top.sv ������һ�� config_db ����
// uvm_config_db#(virtual taxi_axil_if)::set(null, "uvm_test_top.env.slv_agt*", "vif", dut_if);
//         run_test("axil_register_base_test");
//     end

    initial begin
        // Ϊ Master Agent (agt) ���ýӿڣ����������� s_axil (�ӻ���)
        uvm_config_db#(virtual taxi_axil_if)::set(null, "uvm_test_top.env.agt*", "vif", dut_if);
        
        // Ϊ Slave Agent (slv_agt) ���ýӿڣ����������� m_axil (������)
        // ��һ���ǳ��ؼ���Slave Agent �� Driver �������ӵ� Master ��
        uvm_config_db#(virtual taxi_axil_if)::set(null, "uvm_test_top.env.slv_agt*", "vif", dut_if);
        // null�������õ���ʼ·��
        // "uvm_test_top.env.slv_agt*"��Ŀ����������/����·��
        // vif����������ݿ��е�key
        // dut_if����Ҫ���ݵ�ʵ�ʶ�����

        run_test();
    end
endmodule