class axil_register_ral_virt_seq extends axil_register_base_virtual_sequence;
    `uvm_object_utils(axil_register_ral_virt_seq)

    function new(string name = "axil_register_ral_virt_seq");
        super.new(name);
    endfunction

    virtual task body();
        uvm_status_e    status; // ����ʲô��
                                // ����һ��ö�����ͱ��������ڴ�Ų�����ִ�н������ UVM_IS_OK ����ɹ���UVM_NOT_OK ����ʧ�ܣ���ÿ�ε��� read/write ��Ҫ�������
        uvm_reg_data_t  data;   // ������ʲô��
                                // ���� UVM �����һ���������ͣ�Ĭ��ͨ���� 64 λ���߼���������ר��������ŴӼĴ���������д��Ĵ��������ݡ�

        if (rm == null) begin
            `uvm_fatal("RAL_SEQ", "RegModel handle is null!")
        end

        `uvm_info(get_type_name(), "Starting RAL based sequence...", UVM_LOW)

        // --- ���� 1��ǰ��д���� (Frontdoor Write) ---
        // ֱ��ͨ���Ĵ�����дֵ��������״̬���ر�����д������ݣ�·����UVM_FRONTDOOR��
        rm.REG_DATA.write(status, 32'h5555_AAAA, UVM_FRONTDOOR);   // �����write�������ĸ�����ģ�
                                                    // �ú������ն����� uvm_reg �����С���Ϊ��� reg_data �̳��� uvm_reg��������ӵ��������ܡ�
        `uvm_info(get_type_name(), "RAL Write REG_DATA finished", UVM_LOW)

        // --- ���� 2��ǰ�Ŷ����� (Frontdoor Read) ---
        // ������״̬���ر������������ݵĴ�ű�����·��
        rm.REG_DATA.read(status, data);
        `uvm_info(get_type_name(), $sformatf("RAL Read REG_DATA: 'h%0h", data), UVM_LOW)

        // --- ���� 3��ʹ�þ���ֵ�ȶ� ---
        // �������ݺ�RAL ���Զ������ڲ�����ֵ������Լ�鵱ǰӲ��ֵ�Ƿ����Ԥ��
        rm.REG_DATA.mirror(status, UVM_CHECK, UVM_FRONTDOOR);
        
        `uvm_info(get_type_name(), "RAL sequence finished", UVM_LOW)
    endtask
endclass