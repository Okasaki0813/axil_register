class axil_register_write_seq extends uvm_sequence#(axil_register_transaction);
    `uvm_object_utils(axil_register_write_seq)

    // ��������������������� virtual sequence ��ʹ�� with Լ��
    rand bit [31:0] addr;
    rand bit [31:0] data;
    rand bit [3:0]  strb;

    function new(string name = "axil_register_write_seq");
        super.new(name);
    endfunction

    virtual task body();
        // ����һ�� transaction ����

        `uvm_info(get_type_name(), $sformatf("Writing data..."), UVM_LOW)

        req = axil_register_transaction::type_id::create("req");
        
        start_item(req); // ��ʼ����
        
        `uvm_info(get_type_name(), $sformatf("Writing started..."), UVM_LOW)
        
        // �������еı���ֵ���ݸ� transaction
        req.operation = axil_register_transaction::WRITE;
        req.addr      = this.addr;
        req.data      = this.data;
        req.strb      = this.strb;
        
        `uvm_info(get_type_name(), $sformatf("About to finish_item(req) and hand to driver"), UVM_LOW)
        finish_item(req); // �������ֲ����͸� driver

        `uvm_info(get_type_name(), $sformatf("finish_item returned; waiting for driver to complete"), UVM_LOW)

        // ������Եȴ� driver ����Ӧ��ز���ɣ�driver ����� item_done��
        `uvm_info(get_type_name(), $sformatf("Writing data succeed! resp=%0d", req.resp), UVM_LOW)
    endtask
endclass