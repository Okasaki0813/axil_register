`ifndef AXIL_SLAVE_DRIVER_SV
`define AXIL_SLAVE_DRIVER_SV

`include "uvm_macros.svh"

class axil_register_slave_driver extends axil_register_base_driver;
    `uvm_component_utils(axil_register_slave_driver)

    // Slave���е���Ӧ����
    typedef enum {
    RESP_OKAY    = 2'b00,  // �������� OK (Normal Access)
    RESP_EXOKAY  = 2'b01,  // ��ռ���� OK (Exclusive Access OK) - ����ԭ�Ӳ���
    RESP_SLVERR  = 2'b10,  // ���豸���� (Slave Error) - Slave�ڲ�����
    RESP_DECERR  = 2'b11   // ������� (Decode Error) - ��ַ��Ч/δӳ��
} resp_type_t;
    
    resp_type_t default_resp = RESP_OKAY;

    int write_response_delay = 0;
    int read_response_delay = 1;  // ��ͨ��������1�����ӳ�

    // �Ĵ���ģ�ͣ�ģ��Slave�Ĵ洢��
    logic [DATA_W-1:0] register_map [logic [ADDR_W-1:0]];
    
    function new(string name = "axil_slave_driver", uvm_component parent = null);
        super.new(name, parent);
    endfunction

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        
        // ��ȡSlave��������
        if (uvm_config_db#(resp_type_t)::get(this, "", "default_resp", default_resp)) begin
            `uvm_info(get_type_name(), $sformatf("Default response set to %0d", default_resp), UVM_LOW)
        end
    endfunction

    // ����Slave��Ӧ����
    extern task run_phase(uvm_phase phase);

    extern task drive_transaction(axil_register_transaction tr);

    // Slave���з�������Ӧ����ע�⣺��������transaction����
    extern task handle_write_request();
    extern task handle_read_request();

    // ����д��ĸ�������
    extern function void process_write(
        input logic [ADDR_W-1:0] addr,
        input logic [DATA_W-1:0] data,
        input logic [STRB_W-1:0] strb
    );
    
    // �����ȡ�ĸ�������
    extern function void process_read(
        input  logic [ADDR_W-1:0] addr,
        output logic [DATA_W-1:0] data,
        output logic [1:0]        resp
    );
    
    // ��λ���
    extern task wait_for_reset_release();
    
    
endclass

task axil_register_slave_driver::wait_for_reset_release();
    if (vif.rst === 1'b1) begin
        `uvm_info(get_type_name(), "Waiting for reset deassertion", UVM_MEDIUM)
        wait(vif.rst === 1'b0);
        @(posedge vif.clk);
    end
endtask

task axil_register_slave_driver::run_phase(uvm_phase phase);
    // ����slave_driver�е���super.run_phase()����ΪSlave����Ҫ��sequence��ȡtransaction
    
    `uvm_info(get_type_name(), "Slave driver run_phase started", UVM_LOW)
    
    // Slave��������ȡtransaction��������Ӧinterface�ϵ��ź�
    fork
        handle_write_request();  // ��������Ӧд����
        handle_read_request();   // ��������Ӧ������
    join
endtask

task axil_register_slave_driver::drive_transaction(axil_register_transaction tr);
    // Slave driverͨ������Ҫ���������ΪSlave����������transaction
    // ��UVM���Ҫ��ʵ�ִ��麯�������Կ������ջ���Ӿ���
    
    `uvm_info(get_type_name(), 
                 "Slave driver does not actively drive transactions", 
                 UVM_LOW)
endtask

task axil_register_slave_driver::handle_write_request();
    forever begin
        logic [ADDR_W-1:0] awaddr;
        logic [2:0]        awprot;
        logic [DATA_W-1:0] wdata;
        logic [STRB_W-1:0] wstrb;

        // �ȴ�AW��Ч�ź�
        wait(vif.awvalid === 1'b1);
        vif.awready <= 1'b1; // ��ʾ��ģ��׼���ý��յ�ַ

        @(posedge vif.clk iff vif.awvalid && vif.awready);
        awaddr = vif.awaddr;
        awprot = vif.awprot;
        vif.awready <= 1'b0; // ��ַ������ϣ�����ready�ź�

        // �ȴ�W��Ч�ź�
        wait(vif.wvalid === 1'b1);
        vif.wready <= 1'b1; // ��ʾ��ģ��׼���ý�������

        @(posedge vif.clk iff vif.wvalid && vif.wready);
        wdata = vif.wdata;
        wstrb = vif.wstrb;
        vif.wready <= 1'b0; // ���ݽ�����ϣ�����ready�ź�

        `uvm_info(get_type_name(),
                 $sformatf("Received WRITE: addr=0x%0h, data=0x%0h, strb=0x%0h",
                          awaddr, wdata, wstrb),
                 UVM_HIGH)

        // ����д���ӳ�
        repeat(write_response_delay) @(posedge vif.clk);

        // ģ��д��Ĵ���
        process_write(awaddr, wdata, wstrb);

        // ����д��Ӧ
        vif.bresp  <= default_resp;
        vif.bvalid <= 1'b1;

        wait(vif.bready === 1'b1); // �ȴ����豸׼���ý�����Ӧ
        @(posedge vif.clk);
        vif.bvalid <= 1'b0; // ��Ӧ������ϣ�����valid�ź�
    end
endtask

task axil_register_slave_driver::handle_read_request();
    forever begin
        logic [ADDR_W-1:0] araddr;
        logic [2:0]        arprot;

        logic [DATA_W-1:0] rdata;
        logic [1:0]        rresp;

        // �ȴ�AR��Ч�ź�
        wait(vif.arvalid === 1'b1);
        vif.arready <= 1'b1; // ��ʾ��ģ��׼���ý��յ�ַ

        @(posedge vif.clk iff vif.arvalid && vif.arready);
        araddr = vif.araddr;
        arprot = vif.arprot;
        vif.arready <= 1'b0; // ��ַ������ϣ�����ready�ź�

        `uvm_info(get_type_name(),
                 $sformatf("Received READ: addr=0x%0h", araddr),
                 UVM_HIGH)

        // �����ȡ�ӳ�
        repeat(read_response_delay) @(posedge vif.clk);

        // �����ȡ���󣨻�ȡ���ݣ�
        process_read(araddr, rdata, rresp);

        // ���Ͷ���Ӧ
        vif.rdata  <= rdata;
        vif.rresp  <= rresp;
        vif.rvalid <= 1'b1;

        wait(vif.rready === 1'b1); // �ȴ����豸׼���ý�������
        @(posedge vif.clk);
        vif.rvalid <= 1'b0; // ���ݷ�����ϣ�����valid�ź�

        `uvm_info(get_type_name(),
                 $sformatf("Sent READ response: addr=0x%0h, data=0x%0h, resp=%0d",
                          araddr, rdata, rresp),
                 UVM_HIGH)
    end
endtask

function void axil_register_slave_driver::process_write(
    input logic [ADDR_W-1:0] addr,
    input logic [DATA_W-1:0] data,
    input logic [STRB_W-1:0] strb
);
    // ������״η��ʸõ�ַ���ȳ�ʼ��Ϊ0
    if (!register_map.exists(addr)) begin
        register_map[addr] = '0;
    end

    // ����д������¼Ĵ���
    for (int i = 0; i < STRB_W; i++) begin
        if (strb[i]) begin
            register_map[addr][i*8 +: 8] = data[i*8 +: 8];
        end
    end

    `uvm_info(get_type_name(),
             $sformatf("Register at addr=0x%0h updated to 0x%0h",
                      addr, register_map[addr]),
             UVM_HIGH)
endfunction

function void axil_register_slave_driver::process_read(
    input  logic [ADDR_W-1:0] addr,
    output logic [DATA_W-1:0] data,
    output logic [1:0]        resp
);
    // ����ַ�Ƿ���Ч
    if (register_map.exists(addr)) begin
        data = register_map[addr];
        resp = RESP_OKAY;
    end else begin
        // ��ַ��Ч������0�ʹ�����Ӧ
        data = '0;
        resp = RESP_DECERR;  // ��ַ�������
    end
endfunction

`endif // AXIL_REGISTER_SLAVE_DRIVER_SV