`ifndef AXIL_SLAVE_DRIVER_SV
`define AXIL_SLAVE_DRIVER_SV

`include "uvm_macros.svh"

class axil_slave_driver extends axil_register_driver;
    `uvm_component_utils(axil_slave_driver)
    virtual taxi_axil_if vif; // ���鲻Ҫ�ڶ���ʱ�� modport���� connect ʱָ������
    
    // �����༶��ı�־λ�ʹ洢��
    bit aw_done = 1'b0; // д��ַͨ�����ֱ�־λ
    bit w_done  = 1'b0; // д����ͨ�����ֱ�־λ
    logic [31:0] saved_addr; // �����ݴ�awaddr����ֹ2��ʱ�����ں�vif.awaddr�����仯
    bit [31:0] mem_model [bit [31:0]]; // ����������Ϊ Memory Model

    // ��ַ���ƣ�Ĭ��ֵ����������Ĭ����Ϊ��֮ǰһ�£����� 0x0000_3FFF ���� DECERR��
    // ���ǿ����õĳ�Ա��֧��ͨ�� uvm_config_db �� top/test �и��ǡ�
    logic [31:0] addr_limit;

    // RESP ����������ά�����Ķ�
    localparam logic [1:0] RESP_OKAY   = 2'b00;
    localparam logic [1:0] RESP_DECERR = 2'b10;
    function new(string name, uvm_component parent);
        super.new(name, parent);
    endfunction

    // ���� build_phase ����ȡ�ӿ�
    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase); // ������� super��ȷ������� get Ҳ��ִ�У�����еĻ���
        
        // �����ݿ��л�ȡ��Ϊ "vif" �Ľӿڣ�����ֵ�����ص� vif ����
        if (!uvm_config_db#(virtual taxi_axil_if)::get(this, "", "vif", vif)) begin
            `uvm_fatal("SLV_DRV", "Virtual interface not found for slave driver!")
        end

        // ���Դ� config_db ��ȡ��ַ���ޣ����δ������ʹ��Ĭ��ֵ
        if (!uvm_config_db#(logic[31:0])::get(this, "", "addr_limit", addr_limit)) begin
            addr_limit = 32'h0000_3FFF; // backward-compatible default
        end
        `uvm_info(get_type_name(), $sformatf("Slave driver build_phase: vif initialized, addr_limit=0x%0h", addr_limit), UVM_LOW)
    endfunction

    virtual task run_phase(uvm_phase phase);
        int cycle_cnt = 0;

        // ��ʼ����Slave Ĭ������ Ready
        vif.awready <= 1'b1;
        vif.wready  <= 1'b1;
        vif.arready <= 1'b1;
        vif.bvalid  <= 1'b0;
        vif.rvalid  <= 1'b0;

        `uvm_info(get_type_name(), "Slave driver run_phase started", UVM_LOW)

        forever begin
            @(posedge vif.clk);
            if (!vif.rst) begin
                vif.bvalid  <= 1'b0;
                vif.awready <= 1'b1;
                vif.wready  <= 1'b1;
                vif.rvalid  <= 1'b0;
                vif.arready <= 1'b1;
                aw_done     <= 1'b0;
                w_done      <= 1'b0;
                `uvm_info(get_type_name(), "Reset detected, clearing response signals", UVM_LOW)
            end else begin
                // Ĭ�ϱ��� Ready Ϊ 1 (ģ������ӻ�)
                // Ready �ź�Ӧ��Ĭ��Ϊ 1���Ա������ܹ���������
                if (!vif.bvalid) vif.awready <= 1'b1;
                if (!vif.bvalid) vif.wready  <= 1'b1;
                if (!vif.rvalid) vif.arready <= 1'b1;

                // ���������ÿ 200 �Ĵ�ӡһ�ε�ǰ�ź�״̬
                
                cycle_cnt++;
                if ((cycle_cnt % 200) == 0) begin
                    `uvm_info(get_type_name(), $sformatf("Slave running: aw_done=%0b w_done=%0b bvalid=%0b awvalid=%0b awready=%0b wvalid=%0b wready=%0b arready=%0b rvalid=%0b", 
                        aw_done, w_done, vif.bvalid, vif.awvalid, vif.awready, vif.wvalid, vif.wready, vif.arready, vif.rvalid), UVM_MEDIUM)
                end

                // ģ�ⷴѹ��ÿ���� 30% �ĸ������� Ready��ģ��ӻ�æµ
                // vif.awready <= ( $urandom_range(0, 99) < 70 ); 
                // vif.wready  <= ( $urandom_range(0, 99) < 70 );
                // vif.arready <= ( $urandom_range(0, 99) < 70 );
                // `uvm_info("SLV_DRV", $sformatf("awready = 'b%0b, wready = 'b%0b, arready = 'b%0b", vif.awready, vif.wready, vif.arready), UVM_HIGH)
                
                // ע�⣺һ�� valid �� ready ���֣���һ��ͨ��Ҫ�����߼���
                // ����ļ���������ܵ������ֱ���������������Ҫ���Եġ�

                // ������׽��ͨ���������ź�
                if (vif.awvalid && vif.awready) begin 
                    aw_done = 1'b1;
                    saved_addr = vif.awaddr;
                    `uvm_info(get_type_name(), $sformatf("Slave: AW handshake detected, addr=0x%0h", vif.awaddr), UVM_MEDIUM)
                end

                if (vif.wvalid && vif.wready) begin
                    w_done = 1'b1;
                    `uvm_info(get_type_name(), $sformatf("Slave: W handshake detected, data=0x%0h", vif.wdata), UVM_MEDIUM)
                end

                // ����Ƿ�����ͨ�������ֳɹ�����û�н����е�д��Ӧ
                if (aw_done && w_done && !vif.bvalid) begin
                    // �ݴ浱ǰ��������ݣ���ֹ����һ�ĸ���
                    logic [31:0] addr_to_store = saved_addr;
                    logic [31:0] data_to_store = vif.wdata; // ��������ͨ����ʱ�ȶ�
                    logic [31:0] wstrb_mask;    // 32λ����
                    logic [31:0] old_data;      // ԭ������
                    logic [31:0] new_combined_data;

                    `uvm_info(get_type_name(), $sformatf("Slave: Write transaction detected, aw_done=%0b w_done=%0b addr=0x%0h", aw_done, w_done, addr_to_store), UVM_LOW)

                    // �������״̬λ��׼��������һ������ 
                    aw_done = 1'b0; 
                    w_done  = 1'b0;

                    addr_to_store = saved_addr;

                    // ���� 32 λ���룺����λ���Ƽ���
                    // �� wstrb ��ÿһλ��չΪ 8 λ
                    wstrb_mask = {{8{vif.wstrb[3]}}, {8{vif.wstrb[2]}}, {8{vif.wstrb[1]}}, {8{vif.wstrb[0]}}};

                    // ��ȡ�����ݣ������������Ĭ��Ϊ0��
                    old_data = mem_model.exists(addr_to_store) ? mem_model[addr_to_store] : 32'h0;

                    // ������ݣ�(������ & ����) | (������ & ~����)
                    new_combined_data = (vif.wdata & wstrb_mask) | (old_data & ~wstrb_mask);

                    // ���´洢
                    mem_model[addr_to_store] = new_combined_data;

                    `uvm_info("SLV_MEM", $sformatf("WSTRB Write: Addr='h%0h, Data='h%0h, Mask='b%04b, Final='h%0h", 
                    addr_to_store, vif.wdata, vif.wstrb, new_combined_data), UVM_HIGH)

                    fork
                        begin
                            automatic logic [31:0] current_awaddr = saved_addr;
                            `uvm_info(get_type_name(), $sformatf("Slave: B response fork started, will delay 2 cycles then set bvalid, addr=0x%0h", current_awaddr), UVM_LOW)
                            repeat(2) @(posedge vif.clk);   // ģ��ӻ��ӳ�
                                                            // ����ȴ����ܻᵼ��slave�޷���⵽master���͵��µ������źţ��Ӷ�©������
                                                            // ���������ʹ��fork-join_none�ṹ
                            vif.bvalid <= 1'b1;
                            vif.bresp  <= (current_awaddr > addr_limit) ? RESP_DECERR : RESP_OKAY;
                            `uvm_info(get_type_name(), $sformatf("Slave: bvalid set, bresp=0x%0h, waiting for bready...", vif.bresp), UVM_LOW)
                        
                            // ��Ӧ���ֳɹ���Master ���յ� (bready=1)��Slave ���� bvalid
                            do begin
                                @(posedge vif.clk);
                            end while (!vif.bready);

                            vif.bvalid <= 1'b0;
                            `uvm_info(get_type_name(), $sformatf("Slave: bready seen, bvalid cleared, write response complete"), UVM_LOW)
                        end
                    join_none
                end

                if (vif.arvalid && vif.arready && !vif.rvalid) begin
                    `uvm_info("SLV_DRV", $sformatf("Read request received at addr 'h%0h", vif.araddr), UVM_LOW)

                    fork
                        begin
                            automatic logic [31:0] current_araddr = vif.araddr;
                            repeat(2) @(posedge vif.clk);
                            vif.rvalid <= 1'b1;
                            vif.rresp  <= (current_araddr > addr_limit) ? RESP_DECERR : RESP_OKAY;                
                            // --- ��̬��ȡ�洢ģ�� ---
                            if (mem_model.exists(current_araddr)) begin
                                vif.rdata <= mem_model[current_araddr]; // ����֮ǰд����ֵ
                            end else begin
                                vif.rdata <= 32'hDEAD_BEEF; // ���ûд��������һ������ֵ��ʾ��δ���塱
                            end

                            do begin
                                @(posedge vif.clk);
                            end while(!vif.rready);

                            vif.rvalid <= 1'b0;
                        end
                    join_none
                end
            end
        end
    endtask
endclass

`endif // AXIL_SLAVE_DRIVER_SV