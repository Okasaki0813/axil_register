`ifndef AXIL_REGISTER_ADDR_DECODE_VIRT_SEQ_SV
`define AXIL_REGISTER_ADDR_DECODE_VIRT_SEQ_SV

// ��ַ������������ - ���Բ�ͬ��ַ��Χ���ֶ���
class axil_register_addr_decode_virt_seq extends axil_register_base_virtual_sequence;
    `uvm_object_utils(axil_register_addr_decode_virt_seq)

    function new(string name = "axil_register_addr_decode_virt_seq");
        super.new(name);
    endfunction

    virtual task body();
        int test_count = 0;
        int pass_count = 0;

        `uvm_info(get_type_name(), "Starting Address Decode Test...", UVM_LOW)

        // Debug: ��ӡ���� sequencer �е� agt_sqr �Ƿ��ѱ�����
        if (p_sequencer == null) begin
            `uvm_error(get_type_name(), "p_sequencer is null!")
        end else begin
            `uvm_info(get_type_name(), $sformatf("virtual sequencer p_sequencer name = %s", p_sequencer.get_full_name()), UVM_LOW)
            if (p_sequencer.agt_sqr == null) begin
                `uvm_error(get_type_name(), "p_sequencer.agt_sqr is null! Driver sequencer may not be connected.")
            end else begin
                `uvm_info(get_type_name(), $sformatf("agt_sqr name = %s", p_sequencer.agt_sqr.get_full_name()), UVM_LOW)
            end
        end

        // ========== ��һ���֣��Ϸ���ַ��Χ��0x0000_0000 ~ 0x0000_3FFF��- ���� OKAY ==========

        // ���� 1: �����Ϸ���ַд��Ͷ�ȡ����ַ 0��
        test_count++;
        test_write_read_addr_expect_resp(32'h0000_0000, 32'hDEAD_BEEF, 4'hF, 2'b00, pass_count);

        // ���� 2: �Ϸ���Χ�ڵ��м��ַ
        test_count++;
        test_write_read_addr_expect_resp(32'h0000_2000, 32'hCAFE_BABE, 4'hF, 2'b00, pass_count);

        // ���� 3: �Ϸ���Χ�Ͻ磨0x0000_3FFF��
        test_count++;
        test_write_read_addr_expect_resp(32'h0000_3FFC, 32'h1234_5678, 4'hF, 2'b00, pass_count);

        // ���� 4: �Ϸ���Χ�ڵĲ�����д�� - ���ֽ�
        test_count++;
        test_write_read_addr_expect_resp(32'h0000_0004, 32'hXXXX_00FF, 4'b0011, 2'b00, pass_count);

        // ���� 5: �Ϸ���Χ�ڵĲ�����д�� - ���ֽ�
        test_count++;
        test_write_read_addr_expect_resp(32'h0000_0008, 32'hFF00_XXXX, 4'b1100, 2'b00, pass_count);

        // ���� 6: �Ϸ���Χ�ڵ������ַɨ�裨10 �������ַ��
        repeat(10) begin
            bit [31:0] rand_addr;
            bit [31:0] rand_data;
            bit [3:0] rand_strb;
            
            if (!std::randomize(rand_addr) || !std::randomize(rand_data) || !std::randomize(rand_strb)) begin
                `uvm_error(get_type_name(), "Randomization failed")
            end else begin
                // ���������ַ�ںϷ���Χ�ڣ�0x0000_0000 ~ 0x0000_3FFC��
                rand_addr = {14'b0, rand_addr[13:2], 2'b00}; // ��֤�� 0x0~0x3FFC ��Χ�� 4 �ֽڶ���
                test_count++;
                test_write_read_addr_expect_resp(rand_addr, rand_data, rand_strb, 2'b00, pass_count);
            end
        end

        // ========== �ڶ����֣������ַ��Χ��> 0x0000_3FFF��- ���� DECERR ==========

        // ���� 7: �����ַ��0x0000_4000��- Ӧ���� DECERR
        test_count++;
        test_write_read_addr_expect_resp(32'h0000_4000, 32'hBEEF_DEAD, 4'hF, 2'b10, pass_count);

        // ���� 8: ���ߵĳ����ַ��0xFFFF_FFFC��- Ӧ���� DECERR
        test_count++;
        test_write_read_addr_expect_resp(32'hFFFF_FFFC, 32'h9999_8888, 4'hF, 2'b10, pass_count);

        // ���� 9: ��������ַɨ�裨5 ����������ַ��
        repeat(5) begin
            bit [31:0] rand_addr;
            bit [31:0] rand_data;
            bit [3:0] rand_strb;
            
            if (!std::randomize(rand_addr) || !std::randomize(rand_data) || !std::randomize(rand_strb)) begin
                `uvm_error(get_type_name(), "Randomization failed")
            end else begin
                // ���ɳ����ַ���� 0x4000 �� 0xFFFF_FFFC
                // ��֤��ַ��λΪ1��ʹ�� >= 0x4000 �� 4 �ֽڶ���
                rand_addr = {rand_addr[31:15], 1'b1, rand_addr[14:2], 2'b00};
                test_count++;
                test_write_read_addr_expect_resp(rand_addr, rand_data, rand_strb, 2'b10, pass_count);
            end
        end

        // ��ӡ�����ܽ�
        `uvm_info(get_type_name(), $sformatf("Address Decode Test Summary: %0d/%0d tests passed", 
            pass_count, test_count), UVM_LOW)

        if (pass_count == test_count) begin
            `uvm_info(get_type_name(), "All Address Decode Tests PASSED", UVM_LOW)
        end else begin
            `uvm_error(get_type_name(), $sformatf("%0d tests FAILED", test_count - pass_count))
        end
    endtask

    // �������񣺲���д��Ͷ�ȡָ����ַ������֤Ԥ�ڵ���Ӧ��
    virtual task test_write_read_addr_expect_resp(
        bit [31:0] addr, 
        bit [31:0] data, 
        bit [3:0] strb,
        bit [1:0] expected_resp,  // ��������Ӧ�� (OKAY=2'b00 �� DECERR=2'b10)
        output int pass_count     // ���������ͨ���Ĳ�����
    );
    
        axil_register_write_seq wr_seq;
        axil_register_read_seq  rd_seq;
        string resp_name = (expected_resp == 2'b00) ? "OKAY" : "DECERR";

        `uvm_info(get_type_name(), $sformatf("Test: Write to addr 0x%08X, data 0x%08X, strb 4'b%b, expect %s", 
            addr, data, strb, resp_name), UVM_LOW)

        // ִ��д����
        wr_seq = axil_register_write_seq::type_id::create("wr_seq");
        wr_seq.addr = addr;
        wr_seq.data = data;
        wr_seq.strb = strb;
        wr_seq.start(p_sequencer.agt_sqr);  // ֱ���� agt_sqr ����������
        
        // �����Ѿ�������֣����� transaction �а�����Ӧ����
        // ��֤д��Ӧ
        if (wr_seq.req.resp !== expected_resp) begin
            `uvm_error(get_type_name(), $sformatf("Write to addr 0x%08X returned RESP=%0d (expected %s/%02b)", 
                addr, wr_seq.req.resp, resp_name, expected_resp))
        end else begin
            `uvm_info(get_type_name(), $sformatf("Write Response: %s ?", resp_name), UVM_LOW)
            pass_count++;
        end

        // ִ�ж�����
        rd_seq = axil_register_read_seq::type_id::create("rd_seq");
        rd_seq.addr = addr;
        rd_seq.start(p_sequencer.agt_sqr);  // ֱ���� agt_sqr ����������
        
        // �����Ѿ�������֣����� transaction �а�����Ӧ���ݺͶ���������
        // ��֤����Ӧ
        if (rd_seq.req.resp !== expected_resp) begin
            `uvm_error(get_type_name(), $sformatf("Read from addr 0x%08X returned RESP=%0d (expected %s/%02b)", 
                addr, rd_seq.req.resp, resp_name, expected_resp))
        end else begin
            if (expected_resp == 2'b00) begin
                `uvm_info(get_type_name(), $sformatf("Read Response: %s, Data: 0x%08X ?", resp_name, rd_seq.req.data), UVM_LOW)
            end else begin
                `uvm_info(get_type_name(), $sformatf("Read Response: %s ?", resp_name), UVM_LOW)
            end
            pass_count++;
        end
    endtask

endclass

`endif // AXIL_REGISTER_ADDR_DECODE_VIRT_SEQ_SV