`include "uvm_macros.svh"

class axil_register_driver extends uvm_driver#(axil_register_transaction); // #���������driver��Ҫ�����transaction������
    `uvm_component_utils(axil_register_driver)

    virtual taxi_axil_if vif;

    function new(string name = "axil_register_driver", uvm_component parent);
        super.new(name, parent);
    endfunction

    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);
    endfunction

    virtual task run_phase(uvm_phase phase);
        // ��ʼ���źţ���ֹ��ʼ״̬Ϊ����̬
        vif.awvalid <= 0;
        vif.wvalid  <= 0;
        vif.arvalid <= 0;

        forever begin
            seq_item_port.get_next_item(req);
            drive_transfer(req);
            seq_item_port.item_done();
        end
    endtask

    extern task drive_transfer(axil_register_transaction tr);
endclass

task axil_register_driver::drive_transfer(axil_register_transaction tr);
    repeat(tr.delay) @(posedge vif.clk); // Ϊʲô����Ҫ�ȴ�����ʱ�����ڣ�
                                         // ��֤��ͬ�ӳ���ģ�鹤�����ȶ���
                                         // delay�󣬱��ֿ���
                                         // delayС��ʵ����������

    if(tr.operation == axil_register_transaction::WRITE) begin // ΪʲôҪ��WRITEǰ�����axil_register_transaction�����Ӳ�����
                                                               // �ñ������ڱ���WRITE��Ӧ�����������ñ���
        // `uvm_info(get_type_name(), $sformatf("Starting WRITE: addr='h%0h, data='h%0h", tr.addr, tr.data), UVM_LOW)

        fork // �˴�ʹ��fork-join�ṹ��Ϊ��ʵ��д����ͨ����д��ַͨ���ķ��룬��������ͨ����������
            begin // ����AWͨ��
                vif.awaddr  <= tr.addr;
                vif.awprot  <= tr.prot;
                vif.awuser  <= tr.user;
                vif.awvalid <= 1'b1;
                wait(vif.awready == 1'b1);
                @(posedge vif.clk);
                vif.awvalid <= 1'b0;
            end

            begin // ����Wͨ��
                vif.wdata   <= tr.data;
                vif.wstrb   <= tr.strb;
                vif.wuser   <= tr.user;
                vif.wvalid  <= 1'b1;
                wait(vif.wready  == 1'b1);
                @(posedge vif.clk);
                vif.wvalid <= 1'b0;
            end
        join

        vif.bready <= 1'b1; // ��������ģ�飺���Ѿ�׼���ý������д��Ӧ�ź���

        wait(vif.bvalid == 1'b1); // �ȴ�����ģ�����д��Ӧ�ź�

        tr.resp = vif.bresp; // ����Ӧ����������ݰ��У��������scoreboard���м��

        @(posedge vif.clk);
        vif.bready <= 1'b0;

        // `uvm_info(get_type_name(), "AW and W handshake finished.", UVM_HIGH)
    end else if (tr.operation == axil_register_transaction::READ) begin
        vif.araddr  <= tr.addr;
        vif.arprot  <= tr.prot;
        vif.aruser  <= tr.user;
        vif.arvalid <= 1'b1;

        wait(vif.arready == 1'b1);

        @(posedge vif.clk);
        vif.arvalid <= 1'b0;
        vif.rready <= 1'b1;

        wait(vif.rvalid == 1'b1);
        tr.data = vif.rdata;
        tr.resp = vif.rresp;

        // `uvm_info(get_type_name(), $sformatf("Read Back Data: 'h%0h", vif.rdata), UVM_MEDIUM)

        @(posedge vif.clk);
        vif.rready <= 1'b0;
    end
endtask