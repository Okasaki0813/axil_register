`ifndef AXIL_REGISTER_REG_DATA_SV
`define AXIL_REGISTER_REG_DATA_SV

`include "uvm_macros.svh"

class axil_register_reg_data extends uvm_reg;
    `uvm_object_utils(axil_register_reg_data)

    rand uvm_reg_field fld_low;
    rand uvm_reg_field fld_high;

    function new(string name = "axil_register_reg_data");
        // ���������֣���λ���Ƿ�֧�ָ�����
        super.new(name, 32, UVM_NO_COVERAGE);
    endfunction

    virtual function void build();
        fld_low = uvm_reg_field::type_id::create("fld_low");
        fld_low.configure(this, 16, 0, "RW", 0, 16'h0, 1, 1, 1);
        // ������⣺
        // 1. this: ���Ĵ���
        // 2. 16: �ֶ�λ��
        // 3. 0: ���λλ�ã�LSBλ�ã�
        // 4. "RW": ����Ȩ�ޣ�RW/RO/WO�ȣ�
        // 5. 0: �Ƿ���ʧ��volatile����0=����ʧ��1=��ʧ
        // 6. 16'h0: ��λֵ
        // 7. 1: �Ƿ��и�λ��1=�У�
        // 8. 1: �Ƿ���������1=�������
        // 9. 1: �Ƿ�ɵ�����ȡ��1=�ɵ������ʣ�

        fld_high = uvm_reg_field::type_id::create("fld_high");
        // ע�⣺��ʼλ����Ϊ 16
        fld_high.configure(this, 16, 16, "RW", 0, 16'h0, 1, 1, 1);
    endfunction
endclass

`endif // AXIL_REGISTER_REG_DATA_SV